package dutb_scb_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    import dutb_typedef_pkg::*;
    import dutb_util_pkg::*;    
    import dutb_sequence_pkg::*;

    `include "dutb_predictor_base.svh"
    `include "dutb_checker_base.svh"
    `include "dutb_fcc_base.svh"

    `include "dutb_scb_base_cfg.svh"
    `include "dutb_scb_base.svh"
endpackage
