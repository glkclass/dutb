package dutb_macro_pkg;
    `define uvm_debug(a, b) `uvm_info(a, b, UVM_HIGH)
endpackage

