interface dut_if
(
    input clk, rstn
);
endinterface
