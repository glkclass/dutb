/******************************************************************************************************************************
    Project         :   dutb
    Creation Date   :   Dec 2015
    Class           :   dutb_agent_base_cfg
    Description     :   Interface   -   
                        Task        -   
******************************************************************************************************************************/


// ****************************************************************************************************************************
class dutb_agent_base_cfg extends uvm_object;
    `uvm_object_utils(dutb_agent_base_cfg)

    bit                         has_driver, has_monitor;
    dutb_if_proxy_base          dutb_if_h;

    extern function             new(string name = "dutb_agent_base_cfg");
endclass
// ****************************************************************************************************************************


// ****************************************************************************************************************************
function dutb_agent_base_cfg::new(string name = "dutb_agent_base_cfg");
    super.new(name);
    has_driver = 1'b1;
    has_monitor = 1'b1;
endfunction
// ****************************************************************************************************************************



