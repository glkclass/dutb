`timescale 1ns/1ns
package dut_handler_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    import dut_tb_param_pkg::*;
    import typedef_pkg::*;
    `include "dut_handler.svh"
endpackage




