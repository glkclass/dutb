/******************************************************************************************************************************
    Project         :   dutb
    Creation Date   :   Dec 2015
    Class           :   dutb_scb_base_cfg
    Description     :   Interface   -   
                        Task        -   
******************************************************************************************************************************/
// ****************************************************************************************************************************
class dutb_scb_base_cfg extends uvm_object;
    `uvm_object_utils(dutb_scb_base_cfg)

    extern function new(string name = "dutb_scb_base_cfg");
endclass
// ****************************************************************************************************************************


// ****************************************************************************************************************************
function dutb_scb_base_cfg::new(string name = "dutb_scb_base_cfg");
    super.new(name);
endfunction
// ****************************************************************************************************************************



