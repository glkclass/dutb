package dut_env_pkg; 
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    import dut_sequence_pkg::*;
    import dut_agent_pkg::*;
    import dut_scb_pkg::*;
    `include "dut_env_cfg.svh"
    `include "dut_env.svh"
endpackage
