// cpp-class constructor. Creates cpp-class containing all cpp-references(gold references).
import  "DPI-C" function chandle dut_gold_ref_new();

// c-prototype proxy
import  "DPI-C" function void Depth_Rect_dpi
(
    input chandle inst,
    input int in_vec[2 + p_depth_size],
    output int out [p_th_num],
    output int log [p_log_buffer_size]
);


