package dutb_agent_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    import dutb_param_pkg::*;
    import dutb_sequence_pkg::*;
    import dutb_util_pkg::*;
    import dutb_if_proxy_pkg::*;

    `include "dutb_driver_base.svh"
    `include "dutb_monitor_base.svh"
    `include "dutb_agent_base_cfg.svh"
    `include "dutb_agent_base.svh"
endpackage
