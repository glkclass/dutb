package dutb_env_pkg; 
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    import dutb_util_pkg::*;
    import dutb_if_proxy_pkg::*;
    import dutb_sequence_pkg::*;
    import dutb_agent_pkg::*;
    import dutb_scb_pkg::*;
    
    `include "dutb_env_base_cfg.svh"
    `include "dutb_env_base.svh"
endpackage
