`timescale 1ns/1ns

package dutb_util_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    import dutb_param_pkg::*;
    import dutb_typedef_pkg::*;
    import dutb_macro_pkg::*;

    `include "dutb_util.svh"
endpackage

