package dutb_if_proxy_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    `include "dutb_if_proxy_base.svh"
endpackage


 
 
