package dutb_test_pkg;
    `include "uvm_macros.svh"
    import uvm_pkg::*;

    import dutb_typedef_pkg::*;
    import dutb_param_pkg::*;
    import dutb_util_pkg::*;
    import dutb_if_proxy_pkg::*;
    import dutb_env_pkg::*;
    import dutb_agent_pkg::*;
    import dutb_scb_pkg::*;
    import dutb_sequence_pkg::*;
    `include "dutb_test_base.svh"

endpackage




