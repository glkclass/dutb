
interface dutb_if (input clk, rstn);
endinterface
